//module MyInstructionMemory(input logic [7:0]Address,
//						  input clk,
//						  input logic rst,
//						  output logic [15:0]Instruction);
//
//integer i;
//reg [7:0] outputRegister[255:0];
//						  
//always_ff@(posedge clk)
//begin
//
//
//
//	if (RegWr)
//	
//	begin
//	outputRegister[WR] = WD;
//	end
//	
//end
//
//always_comb
//begin
//RD1 = outputRegister[RR1];
//RD2 = outputRegister[RR2];
//end
//
//endmodule

